entity reg4 is 
    port (d0,d1,d2,d3,en,clk) : in bit;
          q0,q1,q2,q3 : out bit );
end entity reg4;

